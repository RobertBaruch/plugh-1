package addr_alu_types;

typedef enum bit[2:0] {
	NONE, INC
} cmd_t /* verilator public */;

endpackage : addr_alu_types
