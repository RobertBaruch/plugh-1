package alu_types;

typedef enum logic[2:0] {
	NONE, OR
} cmd /* verilator public */;

endpackage : alu_types
